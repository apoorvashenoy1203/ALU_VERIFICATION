    package alu_pkg;
  `include "alu_transaction.sv"
  `include "alu_generator.sv"
  `include "alu_driver.sv"
  `include "alu_monitor.sv"
  `include "ref_model.sv"
  `include "scoreboard.sv"
  `include "alu_environment.sv"
  `include "alu_test.sv"
endpackage
